module main

import os
import cli

fn main() {
	println('CLI works!')
}

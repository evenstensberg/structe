module main

fn main() {
	println('CLI works!')
}
